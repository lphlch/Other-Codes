module Divider (
    input I_CLK,
    input rst,
    output O_CLK
);
    
endmodule