`timescale 1ns/1ns
module deselector41_tb;
    reg iS1,iS0,iC;
    reg oZ0,oZ1,oZ2,oZ3;
    deselector41 uut(iC,iS1,iS0,oZ0,oZ1,oZ2,oZ3);
    initial
    begin
        iS1=0;
        iC=0;
        #40 iS1=0;
        #40 iS1=0;
        #40 iS1=1;
        #40 iS1=1;
    end
    initial
    begin
        iS0=0;
        iC=0;
        #40 iS0=0;
        #40 iS0=1;
        #40 iS0=0;
        #40 iS0=1;
    end
endmodule