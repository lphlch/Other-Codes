`timescale 1ns/1ns
module barrelshifter32_tb ();
    reg [31:0] a;
    reg [4:0]  b;
    reg [1:0]  aluc;
    wire [31:0] c;
    barrelshifter32 uut(a,b,aluc,c);
    
    a = 32'b10100101111100001100001111100111;
    
    repeat (31) begin
        b     = 5'b00000;
        #25 b = 5'b00001;
        #25 b = 5'b00010;
        #25 b = 5'b00011;
        #25 b = 5'b00100;
        #25 b = 5'b00101;
        #25 b = 5'b00110;
        #25 b = 5'b00111;
        #25 b = 5'b01000;
        #25 b = 5'b01001;
        #25 b = 5'b01010;
        #25 b = 5'b01011;
        #25 b = 5'b01100;
        #25 b = 5'b01101;
        #25 b = 5'b01110;
        #25 b = 5'b01111;
        #25 b = 5'b10000;
        #25 b = 5'b10001;
        #25 b = 5'b10010;
        #25 b = 5'b10011;
        #25 b = 5'b10100;
        #25 b = 5'b10101;
        #25 b = 5'b10110;
        #25 b = 5'b10111;
        #25 b = 5'b11000;
        #25 b = 5'b11001;
        #25 b = 5'b11010;
        #25 b = 5'b11011;
        #25 b = 5'b11100;
        #25 b = 5'b11101;
        #25 b = 5'b11110;
        #25 b = 5'b11111;
    end
    
    initial begin
        aluc      = 2b'00;
        #800 aluc = 2b'01;
        #800 aluc = 2b'10;
        #800 aluc = 2b'11;
    end
endmodule
